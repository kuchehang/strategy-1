module rconst2in1 (
    i1,
    i2,
    rc1,
    rc2
);
    input [11:0] i1, i2;
    output [63:0] rc1, rc2;
    reg [63:0] rc1, rc2;

    always @(i1) begin
        rc1     = 0;
        rc1[0]  = i1[0] | i1[2] | i1[3] | i1[5] | i1[6] | i1[7] | i1[10] | i1[11];
        rc1[1]  = i1[1] | i1[2] | i1[4] | i1[6] | i1[8] | i1[9];
        rc1[3]  = i1[1] | i1[2] | i1[4] | i1[5] | i1[6] | i1[7] | i1[9];
        rc1[7]  = i1[1] | i1[2] | i1[3] | i1[4] | i1[6] | i1[7] | i1[10];
        rc1[15] = i1[1] | i1[2] | i1[3] | i1[5] | i1[6] | i1[7] | i1[8] | i1[9] | i1[10];
        rc1[31] = i1[3] | i1[5] | i1[6] | i1[10] | i1[11];
        rc1[63] = i1[1] | i1[3] | i1[7] | i1[8] | i1[10];
    end

    always @(i2) begin
        rc2     = 0;
        rc2[0]  = i2[2] | i2[3] | i2[6] | i2[7];
        rc2[1]  = i2[0] | i2[5] | i2[6] | i2[7] | i2[9];
        rc2[3]  = i2[3] | i2[4] | i2[5] | i2[6] | i2[9] | i2[11];
        rc2[7]  = i2[0] | i2[4] | i2[6] | i2[8] | i2[10];
        rc2[15] = i2[0] | i2[1] | i2[3] | i2[7] | i2[10] | i2[11];
        rc2[31] = i2[1] | i2[2] | i2[5] | i2[9] | i2[11];
        rc2[63] = i2[1] | i2[3] | i2[6] | i2[7] | i2[8] | i2[9] | i2[10] | i2[11];
    end
endmodule